** Library name: ECE555_xorcist
** Cell name: OR2
** View name: schematic
mp0 net4 b net1 vdd pmos_rvt w=81e-9 l=20e-9 nfin=3
mp1 net8 a vdd vdd pmos_rvt w=81e-9 l=20e-9 nfin=3
mp2 net4 b net8 vdd pmos_rvt w=81e-9 l=20e-9 nfin=3
mp3 net1 a vdd vdd pmos_rvt w=81e-9 l=20e-9 nfin=3
mp10 y net4 vdd vdd pmos_rvt w=81e-9 l=20e-9 nfin=3
mn4 net4 a vss vss nmos_rvt w=54e-9 l=20e-9 nfin=2
mn0 y net4 vss vss nmos_rvt w=54e-9 l=20e-9 nfin=2
mn5 net4 b vss vss nmos_rvt w=54e-9 l=20e-9 nfin=2
.END
